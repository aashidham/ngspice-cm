* Spice netlister for gnetlist

.control
set temp=300
tran 50us 500ms
plot v(cell_bus) 
.endc



CStray 0 electrode_bus 4e-12
RStray 0 electrode_bus 3e+11
Rbath 0 solution_bus 200.0
Cwholecell solution_bus cell_bus 2e-10
Rwholecell solution_bus cell_bus 100000000.0
R_pene cell_bus Rpene_bus 1e+15
i1 0 cell_bus pulse(0    8e-010      25ms       1ms        1ms        25ms  100ms)
.model memr mig (area=1e-4)
amen cell_bus 0 memr
Xintracpe_i_1 cell_bus electrode_bus cpe_intra_1
Xextracpe_i_1 solution_bus electrode_bus cpe_extra_1

R_seal_i_0 compartment_0 solution_bus 5527741.59845
Xsheathedcpe_i_0 compartment_0 electrode_bus sheathed_cpe_i_0
amen_0 cell_bus compartment_0 memr_0
.model memr_0 trau (area=6.95120334882e-13)
R_seal_i_1 compartment_1 compartment_0 4992923.57323
Xsheathedcpe_i_1 compartment_1 electrode_bus sheathed_cpe_i_1
amen_1 cell_bus compartment_1 memr_1
.model memr_1 trau (area=4.99243932511e-13)
R_seal_i_2 compartment_2 compartment_1 3060019.82182
Xsheathedcpe_i_2 compartment_2 electrode_bus sheathed_cpe_i_2
amen_2 cell_bus compartment_2 memr_2
.model memr_2 trau (area=2.08371941107e-13)
R_seal_i_3 compartment_3 compartment_2 2084171.87382
Xsheathedcpe_i_3 compartment_3 electrode_bus sheathed_cpe_i_3
amen_3 cell_bus compartment_3 memr_3
.model memr_3 trau (area=1.15191730632e-13)
R_seal_i_4 compartment_4 compartment_3 6252515.62147
Xsheathedcpe_i_4 compartment_4 electrode_bus sheathed_cpe_i_4
amen_4 cell_bus compartment_4 memr_4
.model memr_4 trau (area=3.45575191895e-13)
R_seal_i_5 compartment_5 compartment_4 6252515.62147
Xsheathedcpe_i_5 compartment_5 electrode_bus sheathed_cpe_i_5
amen_5 cell_bus compartment_5 memr_5
.model memr_5 trau (area=3.45575191895e-13)
R_seal_i_6 compartment_6 compartment_5 6252515.62147
Xsheathedcpe_i_6 compartment_6 electrode_bus sheathed_cpe_i_6
amen_6 cell_bus compartment_6 memr_6
.model memr_6 trau (area=3.45575191895e-13)
R_seal_i_7 compartment_7 compartment_6 6252515.62147
Xsheathedcpe_i_7 compartment_7 electrode_bus sheathed_cpe_i_7
amen_7 cell_bus compartment_7 memr_7
.model memr_7 trau (area=3.45575191895e-13)

.subckt cpe_intra_1 in out
*k/area=244262588.623 alpha=0.5 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 2.32050730558e+12
c0 rung_0 out 4.30940250692e-07
r1 in rung_1 1.53314397285e+12
c1 rung_1 out 2.84719400115e-07
r2 in rung_2 1.01293817772e+12
c2 rung_2 out 1.88112242177e-07
r3 in rung_3 669241617253.0
c3 rung_3 out 1.24284525896e-07
r4 in rung_4 442163551653.0
c4 rung_4 out 8.21139719483e-08
r5 in rung_5 292134561525.0
c5 rung_5 out 5.42521632561e-08
r6 in rung_6 193011390736.0
c6 rung_6 out 3.58440488035e-08
r7 in rung_7 127521361250.0
c7 rung_7 out 2.36819281946e-08
r8 in rung_8 84252527859.1
c8 rung_8 out 1.56464947943e-08
r9 in rung_9 55665093134.6
c9 rung_9 out 1.03375365949e-08
r10 in rung_10 36777562316.7
c10 rung_10 out 6.82994269679e-09
r11 in rung_11 24298694456.4
c11 rung_11 out 4.51249839004e-09
r12 in rung_12 16053988222.5
c12 rung_12 out 2.98137812044e-09
r13 in rung_13 10606764833.0
c13 rung_13 out 1.96977699021e-09
r14 in rung_14 7007820029.7
c14 rung_14 out 1.30141875147e-09
r15 in rung_15 4630020778.44
c15 rung_15 out 8.59838842209e-10
r16 in rung_16 3059024392.45
c16 rung_16 out 5.6808988939e-10
r17 in rung_17 2021077373.39
c17 rung_17 out 3.75333267799e-10
r18 in rung_18 1335312578.51
c18 rung_18 out 2.47980230854e-10
r19 in rung_19 882232271.667
c19 rung_19 out 1.63838913761e-10
r20 in rung_20 582885081.511
c20 rung_20 out 1.0824729685e-10
r21 in rung_21 385108354.296
c21 rung_21 out 7.15182797936e-11
r22 in rung_22 254438566.456
c22 rung_22 out 4.72516588724e-11
r23 in rung_23 168105893.778
c23 rung_23 out 3.12188614245e-11
r24 in rung_24 111066462.591
c24 rung_24 out 2.06260971974e-11
r25 in rung_25 73380884.127
c25 rung_25 out 1.36275272763e-11
r26 in rung_26 48482269.3517
c26 rung_26 out 9.003617984e-12
r27 in rung_27 32031917.7052
c27 rung_27 out 5.94863141039e-12
r28 in rung_28 21163278.155
c28 rung_28 out 3.93022179746e-12
r29 in rung_29 13982439.2153
c29 rung_29 out 2.5966717908e-12
r30 in rung_30 9238105.97674
c30 rung_30 out 1.71560403881e-12
r31 in rung_31 6103556.09083
c31 rung_31 out 1.13348834781e-12
r32 in rung_32 4032579.51876
c32 rung_32 out 7.48888324794e-13
r33 in rung_33 2664298.86661
c33 rung_33 out 4.94785609481e-13
r34 in rung_34 1760284.80471
c34 rung_34 out 3.26901610352e-13
r35 in rung_35 1163008.6371
c35 rung_35 out 2.15981752103e-13
r36 in rung_36 768392.186506
c36 rung_36 out 1.42697728504e-13
r37 in rung_37 507671.683125
c37 rung_37 out 9.42794542679e-14
r38 in rung_38 335415.35478
c38 rung_38 out 6.22898177165e-14
r39 in rung_39 221606.727264
c39 rung_39 out 4.11544744429e-14
r40 in rung_40 146414.112738
c40 rung_40 out 2.71904916206e-14
r41 in rung_41 96734.8449816
c41 rung_41 out 1.79645796618e-14
r42 in rung_42 63912.0782734
c42 rung_42 out 1.18690800788e-14
r43 in rung_43 42226.2913638
c43 rung_43 out 7.84182344194e-15
r44 in rung_44 27898.6340377
c44 rung_44 out 5.18104136852e-15
r45 in rung_45 18432.4447171
c45 rung_45 out 3.42308008604e-15
r46 in rung_46 12178.1954553
c46 rung_46 out 2.26160658485e-15
r47 in rung_47 8046.0539459
c47 rung_47 out 1.49422865258e-15
r48 in rung_48 5315.97512437
c48 rung_48 out 9.87227080586e-16
r49 in rung_49 3512.22993444
c49 rung_49 out 6.52254463839e-16
rP in out 1.19172262886e+12
cP in out 1.27006168364e-15
.ends

.subckt cpe_extra_1 in out
*k/area=496067355.092 alpha=0.4 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 1.03571616618e+12
c0 rung_0 out 9.65515488369e-07
r1 in rung_1 743431151461.0
c1 rung_1 out 5.87163762754e-07
r2 in rung_2 533630636472.0
c2 rung_2 out 3.57074835613e-07
r3 in rung_3 383037024507.0
c3 rung_3 out 2.17149705612e-07
r4 in rung_4 274941789537.0
c4 rung_4 out 1.320563365e-07
r5 in rung_5 197351646961.0
c5 rung_5 out 8.03080803664e-08
r6 in rung_6 141657885562.0
c6 rung_6 out 4.88381545563e-08
r7 in rung_7 101681221570.0
c7 rung_7 out 2.97001911836e-08
r8 in rung_8 72986200372.3
c8 rung_8 out 1.80617258034e-08
r9 in rung_9 52389077968.9
c9 rung_9 out 1.09839676445e-08
r10 in rung_10 37604581091.0
c10 rung_10 out 6.67973517756e-09
r11 in rung_11 26992353632.8
c11 rung_11 out 4.06218076075e-09
r12 in rung_12 19374957345.6
c12 rung_12 out 2.47035430213e-09
r13 in rung_13 13907233776.3
c13 rung_13 out 1.50230891668e-09
r14 in rung_14 9982533012.0
c14 rung_14 out 9.13606634969e-10
r15 in rung_15 7165405208.44
c15 rung_15 out 5.55596172125e-10
r16 in rung_16 5143286953.26
c16 rung_16 out 3.37877478846e-10
r17 in rung_17 3691822013.42
c17 rung_17 out 2.0547512103e-10
r18 in rung_18 2649968765.62
c18 rung_18 out 1.2495661299e-10
r19 in rung_19 1902132452.01
c19 rung_19 out 7.59904900006e-11
r20 in rung_20 1365339815.3
c20 rung_20 out 4.62124767337e-11
r21 in rung_21 980033125.066
c21 rung_21 out 2.81034245975e-11
r22 in rung_22 703462182.429
c22 rung_22 out 1.70906761536e-11
r23 in rung_23 504941138.673
c23 rung_23 out 1.03934383645e-11
r24 in rung_24 362443866.767
c24 rung_24 out 6.32061365309e-12
r25 in rung_25 260160138.472
c25 rung_25 out 3.843786392e-12
r26 in rung_26 186741462.212
c26 rung_26 out 2.33754104242e-12
r27 in rung_27 134041955.519
c27 rung_27 out 1.42154052482e-12
r28 in rung_28 96214550.4625
c28 rung_28 out 8.64488548878e-13
r29 in rung_29 69062255.0592
c29 rung_29 out 5.25725744778e-13
r30 in rung_30 49572492.4238
c30 rung_30 out 3.19712226473e-13
r31 in rung_31 35582852.0659
c31 rung_31 out 1.94428195255e-13
r32 in rung_32 25541168.0801
c32 rung_32 out 1.1823859077e-13
r33 in rung_33 18333304.6403
c33 rung_33 out 7.1905025549e-14
r34 in rung_34 13159541.4109
c34 rung_34 out 4.37279628042e-14
r35 in rung_35 9445843.70051
c35 rung_35 out 2.65925047158e-14
r36 in rung_36 6780172.68447
c36 rung_36 out 1.61718328894e-14
r37 in rung_37 4866769.24675
c37 rung_37 out 9.83465761486e-15
r38 in rung_38 3493339.18225
c38 rung_38 out 5.98079952119e-15
r39 in rung_39 2507498.92249
c39 rung_39 out 3.63713352447e-15
r40 in rung_40 1799868.41193
c40 rung_40 out 2.21186820055e-15
r41 in rung_41 1291935.27113
c41 rung_41 out 1.34511447097e-15
r42 in rung_42 927343.762307
c42 rung_42 out 8.18011190524e-16
r43 in rung_43 665642.05863
c43 rung_43 out 4.97461236395e-16
r44 in rung_44 477794.069715
c44 rung_44 out 3.02523589631e-16
r45 in rung_45 342957.855644
c45 rung_45 out 1.83975183567e-16
r46 in rung_46 246173.190928
c46 rung_46 out 1.11881748494e-16
r47 in rung_47 176701.711112
c47 rung_47 out 6.80392072634e-17
r48 in rung_48 126835.479494
c48 rung_48 out 4.13770233961e-17
r49 in rung_49 91041.7831117
c49 rung_49 out 2.51628161759e-17
rP in out 407198856654.0
cP in out 3.90501557864e-17
.ends

.subckt sheathed_cpe_i_0 in out
*k/area=431579950.903 alpha=0.5 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 4.10003199696e+12
c0 rung_0 out 2.43900535591e-07
r1 in rung_1 2.70886427701e+12
c1 rung_1 out 1.61143485831e-07
r2 in rung_2 1.78972887936e+12
c2 rung_2 out 1.06466445277e-07
r3 in rung_3 1.18246214431e+12
c3 rung_3 out 7.03416828275e-08
r4 in rung_4 781244991260.0
c4 rung_4 out 4.6474288966e-08
r5 in rung_5 516163447014.0
c5 rung_5 out 3.07052582206e-08
r6 in rung_6 341025807543.0
c6 rung_6 out 2.02867629257e-08
r7 in rung_7 225313516645.0
c7 rung_7 out 1.34033313463e-08
r8 in rung_8 148863164195.0
c8 rung_8 out 8.85549320199e-09
r9 in rung_9 98352917233.4
c9 rung_9 out 5.85076633743e-09
r10 in rung_10 64981128008.5
c10 rung_10 out 3.86556298496e-09
r11 in rung_11 42932605519.4
c11 rung_11 out 2.55395213703e-09
r12 in rung_12 28365291172.5
c12 rung_12 out 1.68737944346e-09
r13 in rung_13 18740762028.5
c13 rung_13 out 1.1148405426e-09
r14 in rung_14 12381898682.9
c14 rung_14 out 7.36567842066e-10
r15 in rung_15 8180639333.7
c15 rung_15 out 4.86645547266e-10
r16 in rung_16 5404894808.29
c16 rung_16 out 3.21523524581e-10
r17 in rung_17 3570978587.01
c17 rung_17 out 2.12428486071e-10
r18 in rung_18 2359322155.41
c18 rung_18 out 1.40350108917e-10
r19 in rung_19 1558788689.82
c19 rung_19 out 9.27283973887e-11
r20 in rung_20 1029881474.19
c20 rung_20 out 6.1265044599e-11
r21 in rung_21 680435942.223
c21 rung_21 out 4.04774135584e-11
r22 in rung_22 449559568.815
c22 rung_22 out 2.67431619304e-11
r23 in rung_23 297021061.606
c23 rung_23 out 1.76690318664e-11
r24 in rung_24 196239869.323
c24 rung_24 out 1.16738135868e-11
r25 in rung_25 129654395.9
c25 rung_25 out 7.71281215004e-12
r26 in rung_26 85661809.8762
c26 rung_26 out 5.09580445324e-12
r27 in rung_27 56596196.5297
c27 rung_27 out 3.36676461459e-12
r28 in rung_28 37392736.2293
c28 rung_28 out 2.22439932184e-12
r29 in rung_29 24705135.8298
c29 rung_29 out 1.46964605769e-12
r30 in rung_30 16322521.3749
c30 rung_30 out 9.70985521208e-13
r31 in rung_31 10784182.9273
c31 rung_31 out 6.41523771972e-13
r32 in rung_32 7125039.00221
c32 rung_32 out 4.23850552883e-13
r33 in rung_33 4707466.58556
c33 rung_33 out 2.80035283224e-13
r34 in rung_34 3110192.3298
c34 rung_34 out 1.85017476837e-13
r35 in rung_35 2054883.69434
c35 rung_35 out 1.22239834713e-13
r36 in rung_36 1357648.19327
c36 rung_36 out 8.07630578806e-14
r37 in rung_37 896989.265991
c37 rung_37 out 5.33596231828e-14
r38 in rung_38 592634.930974
c38 rung_38 out 3.5254353425e-14
r39 in rung_39 391550.015955
c39 rung_39 out 2.32923203216e-14
r40 in rung_40 258694.530109
c40 rung_40 out 1.53890834254e-14
r41 in rung_41 170917.781078
c41 rung_41 out 1.016746659e-14
r42 in rung_42 112924.258106
c42 rung_42 out 6.71757855885e-15
r43 in rung_43 74608.3174519
c43 rung_43 out 4.43826014031e-15
r44 in rung_44 49293.2265074
c44 rung_44 out 2.93232939526e-15
r45 in rung_45 32567.7117846
c45 rung_45 out 1.93737081885e-15
r46 in rung_46 21517.2737927
c46 rung_46 out 1.28000820637e-15
r47 in rung_47 14216.3218138
c47 rung_47 out 8.45693035346e-16
r48 in rung_48 9392.63067715
c48 rung_48 out 5.58743847479e-16
r49 in rung_49 6205.64954795
c49 rung_49 out 3.69158399144e-16
rP in out 2.10561755099e+12
cP in out 7.18820589108e-16
.ends

.subckt sheathed_cpe_i_1 in out
*k/area=600908654.996 alpha=0.5 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 5.70866349926e+12
c0 rung_0 out 1.75172349908e-07
r1 in rung_1 3.77167657084e+12
c1 rung_1 out 1.15735223856e-07
r2 in rung_2 2.49192199836e+12
c2 rung_2 out 7.64655041055e-08
r3 in rung_3 1.64639653726e+12
c3 rung_3 out 5.05202575611e-08
r4 in rung_4 1.08776340499e+12
c4 rung_4 out 3.33784031623e-08
r5 in rung_5 718678154661.0
c5 rung_5 out 2.20528922743e-08
r6 in rung_6 474825948010.0
c6 rung_6 out 1.45702014352e-08
r7 in rung_7 313714392794.0
c7 rung_7 out 9.62643662441e-09
r8 in rung_8 207269043865.0
c8 rung_8 out 6.36012360541e-09
r9 in rung_9 136941299256.0
c9 rung_9 out 4.20209199461e-09
r10 in rung_10 90476219180.4
c10 rung_10 out 2.77629464877e-09
r11 in rung_11 59777045213.0
c11 rung_11 out 1.83427968418e-09
r12 in rung_12 39494302113.5
c12 rung_12 out 1.21189656915e-09
r13 in rung_13 26093626640.0
c13 rung_13 out 8.006921229e-10
r14 in rung_14 17239888155.8
c14 rung_14 out 5.29012039471e-10
r15 in rung_15 11390281148.9
c15 rung_15 out 3.49514788396e-10
r16 in rung_16 7525484126.06
c16 rung_16 out 2.30922130675e-10
r17 in rung_17 4972038055.17
c17 rung_17 out 1.52568738737e-10
r18 in rung_18 3284992966.3
c18 rung_18 out 1.00801166054e-10
r19 in rung_19 2170373329.58
c19 rung_19 out 6.65986699636e-11
r20 in rung_20 1433951438.59
c20 rung_20 out 4.40013048909e-11
r21 in rung_21 947402320.235
c21 rung_21 out 2.90713738452e-11
r22 in rung_22 625942505.606
c22 rung_22 out 1.92072662241e-11
r23 in rung_23 413556112.283
c23 rung_23 out 1.26901149484e-11
r24 in rung_24 273233813.769
c24 rung_24 out 8.38427580088e-12
r25 in rung_25 180523790.531
c25 rung_25 out 5.53943608793e-12
r26 in rung_26 119270885.614
c26 rung_26 out 3.65986912895e-12
r27 in rung_27 78801492.663
c27 rung_27 out 2.41805155406e-12
r28 in rung_28 52063629.8956
c28 rung_28 out 1.59759081872e-12
r29 in rung_29 34398099.1515
c29 rung_29 out 1.05551778652e-12
r30 in rung_30 22726598.7333
c30 rung_30 out 6.97373685811e-13
r31 in rung_31 15015314.8786
c31 rung_31 out 4.60750225028e-13
r32 in rung_32 9920520.16007
c32 rung_32 out 3.04414654844e-13
r33 in rung_33 6554422.67059
c33 rung_33 out 2.01124767933e-13
r34 in rung_34 4330464.11393
c34 rung_34 out 1.32881816405e-13
r35 in rung_35 2861109.26691
c35 rung_35 out 8.77941454584e-14
r36 in rung_36 1890316.14668
c36 rung_36 out 5.80050166778e-14
r37 in rung_37 1248919.49277
c37 rung_37 out 3.83235344706e-14
r38 in rung_38 825152.925964
c38 rung_38 out 2.53201081292e-14
r39 in rung_39 545173.131789
c39 rung_39 out 1.67288295438e-14
r40 in rung_40 360192.316203
c40 rung_40 out 1.10526280724e-14
r41 in rung_41 237976.703338
c41 rung_41 out 7.30239895072e-15
r42 in rung_42 157229.648674
c42 rung_42 out 4.82464714148e-15
r43 in rung_43 103880.598711
c43 rung_43 out 3.18761275532e-15
r44 in rung_44 68633.2309436
c44 rung_44 out 2.10603486223e-15
r45 in rung_45 45345.5260001
c45 rung_45 out 1.39144343475e-15
r46 in rung_46 29959.4919247
c46 rung_46 out 9.19317560612e-16
r47 in rung_47 19794.0400203
c47 rung_47 out 6.07387088935e-16
r48 in rung_48 13077.792551
c48 rung_48 out 4.01296670063e-16
r49 in rung_49 8640.41185285
c49 rung_49 out 2.65134080618e-16
rP in out 2.93174835358e+12
cP in out 5.16265745178e-16
.ends

.subckt sheathed_cpe_i_2 in out
*k/area=1439733192.51 alpha=0.5 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 1.36775402658e+13
c0 rung_0 out 7.31125612183e-08
r1 in rung_1 9.03666123848e+12
c1 rung_1 out 4.8304990164e-08
r2 in rung_2 5.97046287213e+12
c2 rung_2 out 3.19147905074e-08
r3 in rung_3 3.94464570119e+12
c3 rung_3 out 2.10858929828e-08
r4 in rung_4 2.60620156949e+12
c4 rung_4 out 1.39313113391e-08
r5 in rung_5 1.72190030115e+12
c5 rung_5 out 9.20432612391e-09
r6 in rung_6 1.13764824709e+12
c6 rung_6 out 6.08123796339e-09
r7 in rung_7 751636742989.0
c7 rung_7 out 4.01783407819e-09
r8 in rung_8 496601471375.0
c8 rung_8 out 2.65455665064e-09
r9 in rung_9 328101338408.0
c9 rung_9 out 1.75384818644e-09
r10 in rung_10 216774404569.0
c10 rung_10 out 1.15875600558e-09
r11 in rung_11 143221428794.0
c11 rung_11 out 7.65582500728e-10
r12 in rung_12 94625459618.8
c12 rung_12 out 5.05815342141e-10
r13 in rung_13 62518421184.8
c13 rung_13 out 3.34188882454e-10
r14 in rung_14 41305511256.6
c14 rung_14 out 2.20796405034e-10
r15 in rung_15 27290280653.8
c15 rung_15 out 1.4587873815e-10
r16 in rung_16 18030509622.3
c16 rung_16 out 9.63811264992e-11
r17 in rung_17 11912639571.7
c17 rung_17 out 6.36783787896e-11
r18 in rung_18 7870602913.48
c18 rung_18 out 4.2071887646e-11
r19 in rung_19 5200055776.81
c19 rung_19 out 2.77966205131e-11
r20 in rung_20 3435642781.01
c20 rung_20 out 1.83650450497e-11
r21 in rung_21 2269906675.11
c21 rung_21 out 1.21336649367e-11
r22 in rung_22 1499712467.83
c22 rung_22 out 8.01663292401e-12
r23 in rung_23 990850201.392
c23 rung_23 out 5.29653684797e-12
r24 in rung_24 654648236.017
c24 rung_24 out 3.49938719259e-12
r25 in rung_25 432521800.286
c25 rung_25 out 2.31202219018e-12
r26 in rung_26 285764319.569
c26 rung_26 out 1.5275379127e-12
r27 in rung_27 188802613.614
c27 rung_27 out 1.00923429051e-12
r28 in rung_28 124740649.781
c28 rung_28 out 6.66794483242e-13
r29 in rung_29 82415330.0108
c29 rung_29 out 4.40546746246e-13
r30 in rung_30 54451268.5535
c30 rung_30 out 2.91066348786e-13
r31 in rung_31 35975596.369
c31 rung_31 out 1.92305629578e-13
r32 in rung_32 23768840.8092
c32 rung_32 out 1.27055069477e-13
r33 in rung_33 15703917.3894
c33 rung_33 out 8.39444519397e-14
r34 in rung_34 10375475.3272
c34 rung_34 out 5.54615493932e-14
r35 in rung_35 6855008.56864
c35 rung_35 out 3.66430823004e-14
r36 in rung_36 4529059.24734
c36 rung_36 out 2.42098443907e-14
r37 in rung_37 2992319.77036
c37 rung_37 out 1.59952855662e-14
r38 in rung_38 1977006.06662
c38 rung_38 out 1.05679803726e-14
r39 in rung_39 1306194.95489
c39 rung_39 out 6.98219539086e-15
r40 in rung_40 862994.448513
c40 rung_40 out 4.61309074745e-15
r41 in rung_41 570174.7778
c41 rung_41 out 3.0478388319e-15
r42 in rung_42 376710.739911
c42 rung_42 out 2.01368714682e-15
r43 in rung_43 248890.317654
c43 rung_43 out 1.33042990424e-15
r44 in rung_44 164440.202146
c44 rung_44 out 8.79006320766e-16
r45 in rung_45 108644.564147
c45 rung_45 out 5.80753716887e-16
r46 in rung_46 71780.7516936
c46 rung_46 out 3.83700175654e-16
r47 in rung_47 47425.072337
c47 rung_47 out 2.53508192054e-16
r48 in rung_48 31333.4345644
c48 rung_48 out 1.67491201506e-16
r49 in rung_49 20701.7949202
c49 rung_49 out 1.10660339434e-16
rP in out 7.02425465444e+12
cP in out 2.15476420331e-16
.ends

.subckt sheathed_cpe_i_3 in out
*k/area=2604353614.23 alpha=0.5 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 2.47414948897e+13
c0 rung_0 out 4.04179296546e-08
r1 in rung_1 1.63465435675e+13
c1 rung_1 out 2.67038613048e-08
r2 in rung_2 1.08000542326e+13
c2 rung_2 out 1.76430662006e-08
r3 in rung_3 7.13552506962e+12
c3 rung_3 out 1.16566582415e-08
r4 in rung_4 4.71439466159e+12
c4 rung_4 out 7.70147772582e-09
r5 in rung_5 3.11476966424e+12
c5 rung_5 out 5.08831587343e-09
r6 in rung_6 2.05790790921e+12
c6 rung_6 out 3.36181695897e-09
r7 in rung_7 1.35964627222e+12
c7 rung_7 out 2.22113043819e-09
r8 in rung_8 898309383664.0
c8 rung_8 out 1.46748632768e-09
r9 in rung_9 593507124071.0
c9 rung_9 out 9.69558601741e-10
r10 in rung_10 392126268219.0
c10 rung_10 out 6.40581015629e-10
r11 in rung_11 259075256204.0
c11 rung_11 out 4.23227679944e-10
r12 in rung_12 171169324315.0
c12 rung_12 out 2.79623755155e-10
r13 in rung_13 113090451075.0
c13 rung_13 out 1.84745582938e-10
r14 in rung_14 74718120057.4
c14 rung_14 out 1.22060196195e-10
r15 in rung_15 49365772369.3
c15 rung_15 out 8.06443718889e-11
r16 in rung_16 32615642360.3
c16 rung_16 out 5.32812081257e-11
r17 in rung_17 21548941210.0
c17 rung_17 out 3.52025451106e-11
r18 in rung_18 14237244268.9
c18 rung_18 out 2.32580909077e-11
r19 in rung_19 9406454006.17
c19 rung_19 out 1.53664682759e-11
r20 in rung_20 6214782530.86
c20 rung_20 out 1.01525249089e-11
r21 in rung_21 4106066098.93
c21 rung_21 out 6.70770668805e-12
r22 in rung_22 2712850968.65
c22 rung_22 out 4.43173785995e-12
r23 in rung_23 1792362860.41
c23 rung_23 out 2.92802016736e-12
r24 in rung_24 1184202398.32
c24 rung_24 out 1.93452374021e-12
r25 in rung_25 782394765.688
c25 rung_25 out 1.27812716017e-12
r26 in rung_26 516923095.445
c26 rung_26 out 8.44450240445e-13
r27 in rung_27 341527702.284
c27 rung_27 out 5.5792274103e-13
r28 in rung_28 225645115.212
c28 rung_28 out 3.68615899493e-13
r29 in rung_29 149082249.196
c29 rung_29 out 2.43542109627e-13
r30 in rung_30 98497665.2579
c30 rung_30 out 1.60906676144e-13
r31 in rung_31 65076762.0799
c31 rung_31 out 1.06309986669e-13
r32 in rung_32 42995790.3238
c32 rung_32 out 7.02383116501e-14
r33 in rung_33 28407036.9588
c33 rung_33 out 4.64059923063e-14
r34 in rung_34 18768343.196
c34 rung_34 out 3.06601350651e-14
r35 in rung_35 12400121.3796
c35 rung_35 out 2.02569503525e-14
r36 in rung_36 8192678.94997
c36 rung_36 out 1.33836343745e-14
r37 in rung_37 5412849.30388
c37 rung_37 out 8.84247954178e-15
r38 in rung_38 3576234.07012
c38 rung_38 out 5.8421682974e-15
r39 in rung_39 2362794.41867
c39 rung_39 out 3.85988231625e-15
r40 in rung_40 1561082.79141
c40 rung_40 out 2.55019895643e-15
r41 in rung_41 1031397.17208
c41 rung_41 out 1.68489974163e-15
r42 in rung_42 681437.353886
c42 rung_42 out 1.11320221984e-15
r43 in rung_43 450221.19494
c43 rung_43 out 7.35485412957e-16
r44 in rung_44 297458.193651
c44 rung_44 out 4.85930393446e-16
r45 in rung_45 196528.679601
c45 rung_45 out 3.21051027137e-16
r46 in rung_46 129845.210958
c46 rung_46 out 2.12116310106e-16
r47 in rung_47 85787.8801353
c47 rung_47 out 1.40143856302e-16
r48 in rung_48 56679.4903239
c48 rung_48 out 9.25921276376e-17
r49 in rung_49 37447.7678934
c49 rung_49 out 6.11750120672e-17
rP in out 1.27062730037e+13
cP in out 1.19119213635e-16
.ends

.subckt sheathed_cpe_i_4 in out
*k/area=868117871.41 alpha=0.4 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 1.81250329081e+12
c0 rung_0 out 5.51723136211e-07
r1 in rung_1 1.30100451506e+12
c1 rung_1 out 3.35522150145e-07
r2 in rung_2 933853613825.0
c2 rung_2 out 2.04042763208e-07
r3 in rung_3 670314792887.0
c3 rung_3 out 1.24085546064e-07
r4 in rung_4 481148131689.0
c4 rung_4 out 7.54607637144e-08
r5 in rung_5 345365382182.0
c5 rung_5 out 4.58903316379e-08
r6 in rung_6 247901299733.0
c6 rung_6 out 2.79075168893e-08
r7 in rung_7 177942137747.0
c7 rung_7 out 1.69715378192e-08
r8 in rung_8 127725850652.0
c8 rung_8 out 1.03209861734e-08
r9 in rung_9 91680886445.5
c9 rung_9 out 6.27655293974e-09
r10 in rung_10 65808016909.3
c10 rung_10 out 3.81699153003e-09
r11 in rung_11 47236618857.4
c11 rung_11 out 2.321246149e-09
r12 in rung_12 33906175354.8
c12 rung_12 out 1.41163102979e-09
r13 in rung_13 24337659108.5
c13 rung_13 out 8.58462238106e-10
r14 in rung_14 17469432771.0
c14 rung_14 out 5.22060934268e-10
r15 in rung_15 12539459114.8
c15 rung_15 out 3.17483526929e-10
r16 in rung_16 9000752168.21
c16 rung_16 out 1.93072845055e-10
r17 in rung_17 6460688523.49
c17 rung_17 out 1.17414354874e-10
r18 in rung_18 4637445339.84
c18 rung_18 out 7.14037788516e-11
r19 in rung_19 3328731791.02
c19 rung_19 out 4.34231371432e-11
r20 in rung_20 2389344676.77
c20 rung_20 out 2.64071295621e-11
r21 in rung_21 1715057968.86
c21 rung_21 out 1.605909977e-11
r22 in rung_22 1231058819.25
c22 rung_22 out 9.76610065918e-12
r23 in rung_23 883646992.677
c23 rung_23 out 5.93910763686e-12
r24 in rung_24 634276766.843
c24 rung_24 out 3.61177923034e-12
r25 in rung_25 455280242.326
c25 rung_25 out 2.19644936686e-12
r26 in rung_26 326797558.87
c26 rung_26 out 1.33573773852e-12
r27 in rung_27 234573422.158
c27 rung_27 out 8.12308871325e-13
r28 in rung_28 168375463.309
c28 rung_28 out 4.93993456502e-13
r29 in rung_29 120858946.354
c29 rung_29 out 3.00414711301e-13
r30 in rung_30 86751861.7417
c30 rung_30 out 1.82692700841e-13
r31 in rung_31 62269991.1153
c31 rung_31 out 1.1110182586e-13
r32 in rung_32 44697044.1401
c32 rung_32 out 6.75649090113e-14
r33 in rung_33 32083283.1205
c33 rung_33 out 4.1088586028e-14
r34 in rung_34 23029197.4691
c34 rung_34 out 2.49874073167e-14
r35 in rung_35 16530226.4759
c35 rung_35 out 1.51957169805e-14
r36 in rung_36 11865302.1978
c36 rung_36 out 9.24104736536e-15
r37 in rung_37 8516846.1818
c37 rung_37 out 5.61980435135e-15
r38 in rung_38 6113343.56894
c38 rung_38 out 3.41759972639e-15
r39 in rung_39 4388123.11436
c39 rung_39 out 2.07836201398e-15
r40 in rung_40 3149769.72089
c40 rung_40 out 1.26392468603e-15
r41 in rung_41 2260886.72447
c41 rung_41 out 7.68636840555e-16
r42 in rung_42 1622851.58404
c42 rung_42 out 4.67434966014e-16
r43 in rung_43 1164873.6026
c43 rung_43 out 2.84263563654e-16
r44 in rung_44 836139.622
c44 rung_44 out 1.72870622646e-16
r45 in rung_45 600176.247378
c45 rung_45 out 1.05128676324e-16
r46 in rung_46 430803.084124
c46 rung_46 out 6.39324277108e-17
r47 in rung_47 309227.994447
c47 rung_47 out 3.88795470077e-17
r48 in rung_48 221962.089115
c48 rung_48 out 2.36440133692e-17
r49 in rung_49 159323.120445
c49 rung_49 out 1.43787521005e-17
rP in out 712597999144.0
cP in out 2.23143747351e-17
.ends

.subckt sheathed_cpe_i_5 in out
*k/area=868117871.41 alpha=0.4 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 1.81250329081e+12
c0 rung_0 out 5.51723136211e-07
r1 in rung_1 1.30100451506e+12
c1 rung_1 out 3.35522150145e-07
r2 in rung_2 933853613825.0
c2 rung_2 out 2.04042763208e-07
r3 in rung_3 670314792887.0
c3 rung_3 out 1.24085546064e-07
r4 in rung_4 481148131689.0
c4 rung_4 out 7.54607637144e-08
r5 in rung_5 345365382182.0
c5 rung_5 out 4.58903316379e-08
r6 in rung_6 247901299733.0
c6 rung_6 out 2.79075168893e-08
r7 in rung_7 177942137747.0
c7 rung_7 out 1.69715378192e-08
r8 in rung_8 127725850652.0
c8 rung_8 out 1.03209861734e-08
r9 in rung_9 91680886445.5
c9 rung_9 out 6.27655293974e-09
r10 in rung_10 65808016909.3
c10 rung_10 out 3.81699153003e-09
r11 in rung_11 47236618857.4
c11 rung_11 out 2.321246149e-09
r12 in rung_12 33906175354.8
c12 rung_12 out 1.41163102979e-09
r13 in rung_13 24337659108.5
c13 rung_13 out 8.58462238106e-10
r14 in rung_14 17469432771.0
c14 rung_14 out 5.22060934268e-10
r15 in rung_15 12539459114.8
c15 rung_15 out 3.17483526929e-10
r16 in rung_16 9000752168.21
c16 rung_16 out 1.93072845055e-10
r17 in rung_17 6460688523.49
c17 rung_17 out 1.17414354874e-10
r18 in rung_18 4637445339.84
c18 rung_18 out 7.14037788516e-11
r19 in rung_19 3328731791.02
c19 rung_19 out 4.34231371432e-11
r20 in rung_20 2389344676.77
c20 rung_20 out 2.64071295621e-11
r21 in rung_21 1715057968.86
c21 rung_21 out 1.605909977e-11
r22 in rung_22 1231058819.25
c22 rung_22 out 9.76610065918e-12
r23 in rung_23 883646992.677
c23 rung_23 out 5.93910763686e-12
r24 in rung_24 634276766.843
c24 rung_24 out 3.61177923034e-12
r25 in rung_25 455280242.326
c25 rung_25 out 2.19644936686e-12
r26 in rung_26 326797558.87
c26 rung_26 out 1.33573773852e-12
r27 in rung_27 234573422.158
c27 rung_27 out 8.12308871325e-13
r28 in rung_28 168375463.309
c28 rung_28 out 4.93993456502e-13
r29 in rung_29 120858946.354
c29 rung_29 out 3.00414711301e-13
r30 in rung_30 86751861.7417
c30 rung_30 out 1.82692700841e-13
r31 in rung_31 62269991.1153
c31 rung_31 out 1.1110182586e-13
r32 in rung_32 44697044.1401
c32 rung_32 out 6.75649090113e-14
r33 in rung_33 32083283.1205
c33 rung_33 out 4.1088586028e-14
r34 in rung_34 23029197.4691
c34 rung_34 out 2.49874073167e-14
r35 in rung_35 16530226.4759
c35 rung_35 out 1.51957169805e-14
r36 in rung_36 11865302.1978
c36 rung_36 out 9.24104736536e-15
r37 in rung_37 8516846.1818
c37 rung_37 out 5.61980435135e-15
r38 in rung_38 6113343.56894
c38 rung_38 out 3.41759972639e-15
r39 in rung_39 4388123.11436
c39 rung_39 out 2.07836201398e-15
r40 in rung_40 3149769.72089
c40 rung_40 out 1.26392468603e-15
r41 in rung_41 2260886.72447
c41 rung_41 out 7.68636840555e-16
r42 in rung_42 1622851.58404
c42 rung_42 out 4.67434966014e-16
r43 in rung_43 1164873.6026
c43 rung_43 out 2.84263563654e-16
r44 in rung_44 836139.622
c44 rung_44 out 1.72870622646e-16
r45 in rung_45 600176.247378
c45 rung_45 out 1.05128676324e-16
r46 in rung_46 430803.084124
c46 rung_46 out 6.39324277108e-17
r47 in rung_47 309227.994447
c47 rung_47 out 3.88795470077e-17
r48 in rung_48 221962.089115
c48 rung_48 out 2.36440133692e-17
r49 in rung_49 159323.120445
c49 rung_49 out 1.43787521005e-17
rP in out 712597999144.0
cP in out 2.23143747351e-17
.ends

.subckt sheathed_cpe_i_6 in out
*k/area=868117871.41 alpha=0.4 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 1.81250329081e+12
c0 rung_0 out 5.51723136211e-07
r1 in rung_1 1.30100451506e+12
c1 rung_1 out 3.35522150145e-07
r2 in rung_2 933853613825.0
c2 rung_2 out 2.04042763208e-07
r3 in rung_3 670314792887.0
c3 rung_3 out 1.24085546064e-07
r4 in rung_4 481148131689.0
c4 rung_4 out 7.54607637144e-08
r5 in rung_5 345365382182.0
c5 rung_5 out 4.58903316379e-08
r6 in rung_6 247901299733.0
c6 rung_6 out 2.79075168893e-08
r7 in rung_7 177942137747.0
c7 rung_7 out 1.69715378192e-08
r8 in rung_8 127725850652.0
c8 rung_8 out 1.03209861734e-08
r9 in rung_9 91680886445.5
c9 rung_9 out 6.27655293974e-09
r10 in rung_10 65808016909.3
c10 rung_10 out 3.81699153003e-09
r11 in rung_11 47236618857.4
c11 rung_11 out 2.321246149e-09
r12 in rung_12 33906175354.8
c12 rung_12 out 1.41163102979e-09
r13 in rung_13 24337659108.5
c13 rung_13 out 8.58462238106e-10
r14 in rung_14 17469432771.0
c14 rung_14 out 5.22060934268e-10
r15 in rung_15 12539459114.8
c15 rung_15 out 3.17483526929e-10
r16 in rung_16 9000752168.21
c16 rung_16 out 1.93072845055e-10
r17 in rung_17 6460688523.49
c17 rung_17 out 1.17414354874e-10
r18 in rung_18 4637445339.84
c18 rung_18 out 7.14037788516e-11
r19 in rung_19 3328731791.02
c19 rung_19 out 4.34231371432e-11
r20 in rung_20 2389344676.77
c20 rung_20 out 2.64071295621e-11
r21 in rung_21 1715057968.86
c21 rung_21 out 1.605909977e-11
r22 in rung_22 1231058819.25
c22 rung_22 out 9.76610065918e-12
r23 in rung_23 883646992.677
c23 rung_23 out 5.93910763686e-12
r24 in rung_24 634276766.843
c24 rung_24 out 3.61177923034e-12
r25 in rung_25 455280242.326
c25 rung_25 out 2.19644936686e-12
r26 in rung_26 326797558.87
c26 rung_26 out 1.33573773852e-12
r27 in rung_27 234573422.158
c27 rung_27 out 8.12308871325e-13
r28 in rung_28 168375463.309
c28 rung_28 out 4.93993456502e-13
r29 in rung_29 120858946.354
c29 rung_29 out 3.00414711301e-13
r30 in rung_30 86751861.7417
c30 rung_30 out 1.82692700841e-13
r31 in rung_31 62269991.1153
c31 rung_31 out 1.1110182586e-13
r32 in rung_32 44697044.1401
c32 rung_32 out 6.75649090113e-14
r33 in rung_33 32083283.1205
c33 rung_33 out 4.1088586028e-14
r34 in rung_34 23029197.4691
c34 rung_34 out 2.49874073167e-14
r35 in rung_35 16530226.4759
c35 rung_35 out 1.51957169805e-14
r36 in rung_36 11865302.1978
c36 rung_36 out 9.24104736536e-15
r37 in rung_37 8516846.1818
c37 rung_37 out 5.61980435135e-15
r38 in rung_38 6113343.56894
c38 rung_38 out 3.41759972639e-15
r39 in rung_39 4388123.11436
c39 rung_39 out 2.07836201398e-15
r40 in rung_40 3149769.72089
c40 rung_40 out 1.26392468603e-15
r41 in rung_41 2260886.72447
c41 rung_41 out 7.68636840555e-16
r42 in rung_42 1622851.58404
c42 rung_42 out 4.67434966014e-16
r43 in rung_43 1164873.6026
c43 rung_43 out 2.84263563654e-16
r44 in rung_44 836139.622
c44 rung_44 out 1.72870622646e-16
r45 in rung_45 600176.247378
c45 rung_45 out 1.05128676324e-16
r46 in rung_46 430803.084124
c46 rung_46 out 6.39324277108e-17
r47 in rung_47 309227.994447
c47 rung_47 out 3.88795470077e-17
r48 in rung_48 221962.089115
c48 rung_48 out 2.36440133692e-17
r49 in rung_49 159323.120445
c49 rung_49 out 1.43787521005e-17
rP in out 712597999144.0
cP in out 2.23143747351e-17
.ends

.subckt sheathed_cpe_i_7 in out
*k/area=868117871.41 alpha=0.4 n=50 f_low=1e-06 f_high=1e+12
r0 in rung_0 1.81250329081e+12
c0 rung_0 out 5.51723136211e-07
r1 in rung_1 1.30100451506e+12
c1 rung_1 out 3.35522150145e-07
r2 in rung_2 933853613825.0
c2 rung_2 out 2.04042763208e-07
r3 in rung_3 670314792887.0
c3 rung_3 out 1.24085546064e-07
r4 in rung_4 481148131689.0
c4 rung_4 out 7.54607637144e-08
r5 in rung_5 345365382182.0
c5 rung_5 out 4.58903316379e-08
r6 in rung_6 247901299733.0
c6 rung_6 out 2.79075168893e-08
r7 in rung_7 177942137747.0
c7 rung_7 out 1.69715378192e-08
r8 in rung_8 127725850652.0
c8 rung_8 out 1.03209861734e-08
r9 in rung_9 91680886445.5
c9 rung_9 out 6.27655293974e-09
r10 in rung_10 65808016909.3
c10 rung_10 out 3.81699153003e-09
r11 in rung_11 47236618857.4
c11 rung_11 out 2.321246149e-09
r12 in rung_12 33906175354.8
c12 rung_12 out 1.41163102979e-09
r13 in rung_13 24337659108.5
c13 rung_13 out 8.58462238106e-10
r14 in rung_14 17469432771.0
c14 rung_14 out 5.22060934268e-10
r15 in rung_15 12539459114.8
c15 rung_15 out 3.17483526929e-10
r16 in rung_16 9000752168.21
c16 rung_16 out 1.93072845055e-10
r17 in rung_17 6460688523.49
c17 rung_17 out 1.17414354874e-10
r18 in rung_18 4637445339.84
c18 rung_18 out 7.14037788516e-11
r19 in rung_19 3328731791.02
c19 rung_19 out 4.34231371432e-11
r20 in rung_20 2389344676.77
c20 rung_20 out 2.64071295621e-11
r21 in rung_21 1715057968.86
c21 rung_21 out 1.605909977e-11
r22 in rung_22 1231058819.25
c22 rung_22 out 9.76610065918e-12
r23 in rung_23 883646992.677
c23 rung_23 out 5.93910763686e-12
r24 in rung_24 634276766.843
c24 rung_24 out 3.61177923034e-12
r25 in rung_25 455280242.326
c25 rung_25 out 2.19644936686e-12
r26 in rung_26 326797558.87
c26 rung_26 out 1.33573773852e-12
r27 in rung_27 234573422.158
c27 rung_27 out 8.12308871325e-13
r28 in rung_28 168375463.309
c28 rung_28 out 4.93993456502e-13
r29 in rung_29 120858946.354
c29 rung_29 out 3.00414711301e-13
r30 in rung_30 86751861.7417
c30 rung_30 out 1.82692700841e-13
r31 in rung_31 62269991.1153
c31 rung_31 out 1.1110182586e-13
r32 in rung_32 44697044.1401
c32 rung_32 out 6.75649090113e-14
r33 in rung_33 32083283.1205
c33 rung_33 out 4.1088586028e-14
r34 in rung_34 23029197.4691
c34 rung_34 out 2.49874073167e-14
r35 in rung_35 16530226.4759
c35 rung_35 out 1.51957169805e-14
r36 in rung_36 11865302.1978
c36 rung_36 out 9.24104736536e-15
r37 in rung_37 8516846.1818
c37 rung_37 out 5.61980435135e-15
r38 in rung_38 6113343.56894
c38 rung_38 out 3.41759972639e-15
r39 in rung_39 4388123.11436
c39 rung_39 out 2.07836201398e-15
r40 in rung_40 3149769.72089
c40 rung_40 out 1.26392468603e-15
r41 in rung_41 2260886.72447
c41 rung_41 out 7.68636840555e-16
r42 in rung_42 1622851.58404
c42 rung_42 out 4.67434966014e-16
r43 in rung_43 1164873.6026
c43 rung_43 out 2.84263563654e-16
r44 in rung_44 836139.622
c44 rung_44 out 1.72870622646e-16
r45 in rung_45 600176.247378
c45 rung_45 out 1.05128676324e-16
r46 in rung_46 430803.084124
c46 rung_46 out 6.39324277108e-17
r47 in rung_47 309227.994447
c47 rung_47 out 3.88795470077e-17
r48 in rung_48 221962.089115
c48 rung_48 out 2.36440133692e-17
r49 in rung_49 159323.120445
c49 rung_49 out 1.43787521005e-17
rP in out 712597999144.0
cP in out 2.23143747351e-17
.ends
